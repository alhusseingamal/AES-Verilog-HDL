module InvSBox(xy, xy_out);
    
    input [7:0] xy;
    output reg [7:0] xy_out;

    always @(xy) begin  
        case(xy)
            8'h00: xy_out = 8'h52;
            8'h01: xy_out = 8'h09;
            8'h02: xy_out = 8'h6a;
            8'h03: xy_out = 8'hd5;
            8'h04: xy_out = 8'h30;
            8'h05: xy_out = 8'h36;
            8'h06: xy_out = 8'ha5;
            8'h07: xy_out = 8'h38;
            8'h08: xy_out = 8'hbf;
            8'h09: xy_out = 8'h40;
            8'h0a: xy_out = 8'ha3;
            8'h0b: xy_out = 8'h9e;
            8'h0c: xy_out = 8'h81;
            8'h0d: xy_out = 8'hf3;
            8'h0e: xy_out = 8'hd7;
            8'h0f: xy_out = 8'hfb;
            8'h10: xy_out = 8'h7c;
            8'h11: xy_out = 8'he3;
            8'h12: xy_out = 8'h39;
            8'h13: xy_out = 8'h82;
            8'h14: xy_out = 8'h9b;
            8'h15: xy_out = 8'h2f;
            8'h16: xy_out = 8'hff;
            8'h17: xy_out = 8'h87;
            8'h18: xy_out = 8'h34;
            8'h19: xy_out = 8'h8e;
            8'h1a: xy_out = 8'h43;
            8'h1b: xy_out = 8'h44;
            8'h1c: xy_out = 8'hc4;
            8'h1d: xy_out = 8'hde;
            8'h1e: xy_out = 8'he9;
            8'h1f: xy_out = 8'hcb;
            8'h20: xy_out = 8'h54;
            8'h21: xy_out = 8'h7b;
            8'h22: xy_out = 8'h94;
            8'h23: xy_out = 8'h32;
            8'h24: xy_out = 8'ha6;
            8'h25: xy_out = 8'hc2;
            8'h26: xy_out = 8'h23;
            8'h27: xy_out = 8'h3d;
            8'h28: xy_out = 8'hee;
            8'h29: xy_out = 8'h4c;
            8'h2a: xy_out = 8'h95;
            8'h2b: xy_out = 8'h0b;
            8'h2c: xy_out = 8'h42;
            8'h2d: xy_out = 8'hfa;
            8'h2e: xy_out = 8'hc3;
            8'h2f: xy_out = 8'h4e;
            8'h30: xy_out = 8'h08;
            8'h31: xy_out = 8'h2e;
            8'h32: xy_out = 8'ha1;
            8'h33: xy_out = 8'h66;
            8'h34: xy_out = 8'h28;
            8'h35: xy_out = 8'hd9;
            8'h36: xy_out = 8'h24;
            8'h37: xy_out = 8'hb2;
            8'h38: xy_out = 8'h76;
            8'h39: xy_out = 8'h5b;
            8'h3a: xy_out = 8'ha2;
            8'h3b: xy_out = 8'h49;
            8'h3c: xy_out = 8'h6d;
            8'h3d: xy_out = 8'h8b;
            8'h3e: xy_out = 8'hd1;
            8'h3f: xy_out = 8'h25;
            8'h40: xy_out = 8'h72;
            8'h41: xy_out = 8'hf8;
            8'h42: xy_out = 8'hf6;
            8'h43: xy_out = 8'h64;
            8'h44: xy_out = 8'h86;
            8'h45: xy_out = 8'h68;
            8'h46: xy_out = 8'h98;
            8'h47: xy_out = 8'h16;
            8'h48: xy_out = 8'hd4;
            8'h49: xy_out = 8'ha4;
            8'h4a: xy_out = 8'h5c;
            8'h4b: xy_out = 8'hcc;
            8'h4c: xy_out = 8'h5d;
            8'h4d: xy_out = 8'h65;
            8'h4e: xy_out = 8'hb6;
            8'h4f: xy_out = 8'h92;
            8'h50: xy_out = 8'h6c;
            8'h51: xy_out = 8'h70;
            8'h52: xy_out = 8'h48;
            8'h53: xy_out = 8'h50;
            8'h54: xy_out = 8'hfd;
            8'h55: xy_out = 8'hed;
            8'h56: xy_out = 8'hb9;
            8'h57: xy_out = 8'hda;
            8'h58: xy_out = 8'h5e;
            8'h59: xy_out = 8'h15;
            8'h5a: xy_out = 8'h46;
            8'h5b: xy_out = 8'h57;
            8'h5c: xy_out = 8'ha7;
            8'h5d: xy_out = 8'h8d;
            8'h5e: xy_out = 8'h9d;
            8'h5f: xy_out = 8'h84;
            8'h60: xy_out = 8'h90;
            8'h61: xy_out = 8'hd8;
            8'h62: xy_out = 8'hab;
            8'h63: xy_out = 8'h00;
            8'h64: xy_out = 8'h8c;
            8'h65: xy_out = 8'hbc;
            8'h66: xy_out = 8'hd3;
            8'h67: xy_out = 8'h0a;
            8'h68: xy_out = 8'hf7;
            8'h69: xy_out = 8'he4;
            8'h6a: xy_out = 8'h58;
            8'h6b: xy_out = 8'h05;
            8'h6c: xy_out = 8'hb8;
            8'h6d: xy_out = 8'hb3;
            8'h6e: xy_out = 8'h45;
            8'h6f: xy_out = 8'h06;
            8'h70: xy_out = 8'hd0;
            8'h71: xy_out = 8'h2c;
            8'h72: xy_out = 8'h1e;
            8'h73: xy_out = 8'h8f;
            8'h74: xy_out = 8'hca;
            8'h75: xy_out = 8'h3f;
            8'h76: xy_out = 8'h0f;
            8'h77: xy_out = 8'h02;
            8'h78: xy_out = 8'hc1;
            8'h79: xy_out = 8'haf;
            8'h7a: xy_out = 8'hbd;
            8'h7b: xy_out = 8'h03;
            8'h7c: xy_out = 8'h01;
            8'h7d: xy_out = 8'h13;
            8'h7e: xy_out = 8'h8a;
            8'h7f: xy_out = 8'h6b;
            8'h80: xy_out = 8'h3a;
            8'h81: xy_out = 8'h91;
            8'h82: xy_out = 8'h11;
            8'h83: xy_out = 8'h41;
            8'h84: xy_out = 8'h4f;
            8'h85: xy_out = 8'h67;
            8'h86: xy_out = 8'hdc;
            8'h87: xy_out = 8'hea;
            8'h88: xy_out = 8'h97;
            8'h89: xy_out = 8'hf2;
            8'h8a: xy_out = 8'hcf;
            8'h8b: xy_out = 8'hce;
            8'h8c: xy_out = 8'hf0;
            8'h8d: xy_out = 8'hb4;
            8'h8e: xy_out = 8'he6;
            8'h8f: xy_out = 8'h73;
            8'h90: xy_out = 8'h96;
            8'h91: xy_out = 8'hac;
            8'h92: xy_out = 8'h74;
            8'h93: xy_out = 8'h22;
            8'h94: xy_out = 8'he7;
            8'h95: xy_out = 8'had;
            8'h96: xy_out = 8'h35;
            8'h97: xy_out = 8'h85;
            8'h98: xy_out = 8'he2;
            8'h99: xy_out = 8'hf9;
            8'h9a: xy_out = 8'h37;
            8'h9b: xy_out = 8'he8;
            8'h9c: xy_out = 8'h1c;
            8'h9d: xy_out = 8'h75;
            8'h9e: xy_out = 8'hdf;
            8'h9f: xy_out = 8'h6e;
            8'ha0: xy_out = 8'h47;
            8'ha1: xy_out = 8'hf1;
            8'ha2: xy_out = 8'h1a;
            8'ha3: xy_out = 8'h71;
            8'ha4: xy_out = 8'h1d;
            8'ha5: xy_out = 8'h29;
            8'ha6: xy_out = 8'hc5;
            8'ha7: xy_out = 8'h89;
            8'ha8: xy_out = 8'h6f;
            8'ha9: xy_out = 8'hb7;
            8'haa: xy_out = 8'h62;
            8'hab: xy_out = 8'h0e;
            8'hac: xy_out = 8'haa;
            8'had: xy_out = 8'h18;
            8'hae: xy_out = 8'hbe;
            8'haf: xy_out = 8'h1b;
            8'hb0: xy_out = 8'hfc;
            8'hb1: xy_out = 8'h56;
            8'hb2: xy_out = 8'h3e;
            8'hb3: xy_out = 8'h4b;
            8'hb4: xy_out = 8'hc6;
            8'hb5: xy_out = 8'hd2;
            8'hb6: xy_out = 8'h79;
            8'hb7: xy_out = 8'h20;
            8'hb8: xy_out = 8'h9a;
            8'hb9: xy_out = 8'hdb;
            8'hba: xy_out = 8'hc0;
            8'hbb: xy_out = 8'hfe;
            8'hbc: xy_out = 8'h78;
            8'hbd: xy_out = 8'hcd;
            8'hbe: xy_out = 8'h5a;
            8'hbf: xy_out = 8'hf4;
            8'hc0: xy_out = 8'h1f;
            8'hc1: xy_out = 8'hdd;
            8'hc2: xy_out = 8'ha8;
            8'hc3: xy_out = 8'h33;
            8'hc4: xy_out = 8'h88;
            8'hc5: xy_out = 8'h07;
            8'hc6: xy_out = 8'hc7;
            8'hc7: xy_out = 8'h31;
            8'hc8: xy_out = 8'hb1;
            8'hc9: xy_out = 8'h12;
            8'hca: xy_out = 8'h10;
            8'hcb: xy_out = 8'h59;
            8'hcc: xy_out = 8'h27;
            8'hcd: xy_out = 8'h80;
            8'hce: xy_out = 8'hec;
            8'hcf: xy_out = 8'h5f;
            8'hd0: xy_out = 8'h60;
            8'hd1: xy_out = 8'h51;
            8'hd2: xy_out = 8'h7f;
            8'hd3: xy_out = 8'ha9;
            8'hd4: xy_out = 8'h19;
            8'hd5: xy_out = 8'hb5;
            8'hd6: xy_out = 8'h4a;
            8'hd7: xy_out = 8'h0d;
            8'hd8: xy_out = 8'h2d;
            8'hd9: xy_out = 8'he5;
            8'hda: xy_out = 8'h7a;
            8'hdb: xy_out = 8'h9f;
            8'hdc: xy_out = 8'h93;
            8'hdd: xy_out = 8'hc9;
            8'hde: xy_out = 8'h9c;
            8'hdf: xy_out = 8'hef;
            8'he0: xy_out = 8'ha0;
            8'he1: xy_out = 8'he0;
            8'he2: xy_out = 8'h3b;
            8'he3: xy_out = 8'h4d;
            8'he4: xy_out = 8'hae;
            8'he5: xy_out = 8'h2a;
            8'he6: xy_out = 8'hf5;
            8'he7: xy_out = 8'hb0;
            8'he8: xy_out = 8'hc8;
            8'he9: xy_out = 8'heb;
            8'hea: xy_out = 8'hbb;
            8'heb: xy_out = 8'h3c;
            8'hec: xy_out = 8'h83;
            8'hed: xy_out = 8'h53;
            8'hee: xy_out = 8'h99;
            8'hef: xy_out = 8'h61;
            8'hf0: xy_out = 8'h17;
            8'hf1: xy_out = 8'h2b;
            8'hf2: xy_out = 8'h04;
            8'hf3: xy_out = 8'h7e;
            8'hf4: xy_out = 8'hba;
            8'hf5: xy_out = 8'h77;
            8'hf6: xy_out = 8'hd6;
            8'hf7: xy_out = 8'h26;
            8'hf8: xy_out = 8'he1;
            8'hf9: xy_out = 8'h69;
            8'hfa: xy_out = 8'h14;
            8'hfb: xy_out = 8'h63;
            8'hfc: xy_out = 8'h55;
            8'hfd: xy_out = 8'h21;
            8'hfe: xy_out = 8'h0c;
            8'hff: xy_out = 8'h7d;
        endcase
    end
endmodule